
`define data_width 8